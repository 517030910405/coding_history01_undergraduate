module mem_reader(
	input wire [63:0] clk_cnt;
	input wire enable;
	output wire ready;
	input wire w;
	input wire [31:0] addr;
	input wire [7:0] data_in;
	output wire [7:0] data_out;
);
	always @(clk_cnt or ) begin
		
		
		
	end
	
	
endmodule